interface idu_exu_if (
    input logic clk
);
  logic [ 3:0] rd;
  logic [31:0] imm;
endinterface
