`include "ysyx_macro.svh"
