`include "ysyx_macro.vh"
