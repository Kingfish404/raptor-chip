// 触发器模板
module ysyx_Reg (
  input clk,
  input rst,
  input [WIDTH-1:0] din,
  output reg [WIDTH-1:0] dout,
  input wen
);
  parameter WIDTH = 1;
  parameter RESET_VAL = 0;
  always @(posedge clk) begin
    if (rst) dout <= RESET_VAL;
    else if (wen) dout <= din;
  end
endmodule

// // 使用触发器模板的示例
// module example(
//   input clk,
//   input rst,
//   input [3:0] in,
//   output [3:0] out
// );
//   // 位宽为1比特, 复位值为1'b1, 写使能一直有效
//   Reg #(1, 1'b1) i0 (clk, rst, in[0], out[0], 1'b1);
//   // 位宽为3比特, 复位值为3'b0, 写使能为out[0]
//   Reg #(3, 3'b0) i1 (clk, rst, in[3:1], out[3:1], out[0]);
// endmodule

// // 选择器模板内部实现
// module MuxKeyInternal (
//   output reg [DATA_LEN-1:0] out,
//   input [KEY_LEN-1:0] key,
//   input [DATA_LEN-1:0] default_out,
//   input [NR_KEY*(KEY_LEN + DATA_LEN)-1:0] lut
// );
//   parameter NR_KEY = 2;
//   parameter KEY_LEN = 1;
//   parameter DATA_LEN = 1;
//   parameter HAS_DEFAULT = 0;

//   localparam PAIR_LEN = KEY_LEN + DATA_LEN;
//   wire [PAIR_LEN-1:0] pair_list [NR_KEY-1:0];
//   wire [KEY_LEN-1:0] key_list [NR_KEY-1:0];
//   wire [DATA_LEN-1:0] data_list [NR_KEY-1:0];

//   generate
//     for (genvar n = 0; n < NR_KEY; n = n + 1) begin
//       assign pair_list[n] = lut[PAIR_LEN*(n+1)-1 : PAIR_LEN*n];
//       assign data_list[n] = pair_list[n][DATA_LEN-1:0];
//       assign key_list[n]  = pair_list[n][PAIR_LEN-1:DATA_LEN];
//     end
//   endgenerate

//   reg [DATA_LEN-1 : 0] lut_out;
//   reg hit;
//   integer i;
//   always @(*) begin
//     lut_out = 0;
//     hit = 0;
//     for (i = 0; i < NR_KEY; i = i + 1) begin
//       lut_out = lut_out | ({DATA_LEN{key == key_list[i]}} & data_list[i]);
//       hit = hit | (key == key_list[i]);
//     end
//     if (!HAS_DEFAULT) out = lut_out;
//     else out = (hit ? lut_out : default_out);
//   end
// endmodule

// // 不带默认值的选择器模板
// module MuxKey (
//   output [DATA_LEN-1:0] out,
//   input [KEY_LEN-1:0] key,
//   input [NR_KEY*(KEY_LEN + DATA_LEN)-1:0] lut
// );
//   parameter NR_KEY = 2;
//   parameter KEY_LEN = 1;
//   parameter DATA_LEN = 1;
//   MuxKeyInternal #(NR_KEY, KEY_LEN, DATA_LEN, 0) i0 (out, key, {DATA_LEN{1'b0}}, lut);
// endmodule

// // 带默认值的选择器模板
// module MuxKeyWithDefault (
//   output [DATA_LEN-1:0] out,
//   input [KEY_LEN-1:0] key,
//   input [DATA_LEN-1:0] default_out,
//   input [NR_KEY*(KEY_LEN + DATA_LEN)-1:0] lut
// );
//   parameter NR_KEY = 2;
//   parameter KEY_LEN = 1;
//   parameter DATA_LEN = 1;
//   MuxKeyInternal #(NR_KEY, KEY_LEN, DATA_LEN, 1) i0 (out, key, default_out, lut);
// endmodule


// // 使用选择器模板来分别实现2选1多路选择器和4选1多路选择器:
// module mux21(a,b,s,y);
//   input   a,b,s;
//   output  y;

//   // 通过MuxKey实现如下always代码
//   // always @(*) begin
//   //  case (s)
//   //    1'b0: y = a;
//   //    1'b1: y = b;
//   //  endcase
//   // end
//   MuxKey #(2, 1, 1) i0 (y, s, {
//     1'b0, a,
//     1'b1, b
//   });
// endmodule

// module mux41(a,s,y);
//   input  [3:0] a;
//   input  [1:0] s;
//   output y;

//   // 通过MuxKeyWithDefault实现如下always代码
//   // always @(*) begin
//   //  case (s)
//   //    2'b00: y = a[0];
//   //    2'b01: y = a[1];
//   //    2'b10: y = a[2];
//   //    2'b11: y = a[3];
//   //    default: y = 1'b0;
//   //  endcase
//   // end
//   MuxKeyWithDefault #(4, 2, 1) i0 (y, s, 1'b0, {
//     2'b00, a[0],
//     2'b01, a[1],
//     2'b10, a[2],
//     2'b11, a[3]
//   });
// endmodule