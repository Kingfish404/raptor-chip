`include "ysyx.svh"
